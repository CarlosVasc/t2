
.options savecurrents

.include ../doc/ngspice_5.txt

.control

*makes plots in color
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0

echo "********************************************"
echo  "Transient analysis"
echo "********************************************"
tran 1e-6 20e-3 uic



hardcopy Simulacao4.eps v(V6) v(V1) 


quit

.endc
.end
